module system(input a, output b);

	assign b = !a;

endmodule

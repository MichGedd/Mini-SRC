module shift_mask_32 (input [4:0] in_shift, input in_left, output reg [31:0] out_mask);
	
	// in_left = 1 -> shift/rot left
	// in_left = 0 -> shift/rot right
	
	always @(*) begin
		case(in_left)
			1'b0 : begin  // shift right
				case(in_shift)
					5'b00000: out_mask = 32'b11111111111111111111111111111111;
					5'b00001: out_mask = 32'b1111111111111111111111111111111;
					5'b00010: out_mask = 32'b111111111111111111111111111111;
					5'b00011: out_mask = 32'b11111111111111111111111111111;
					5'b00100: out_mask = 32'b1111111111111111111111111111;
					5'b00101: out_mask = 32'b111111111111111111111111111;
					5'b00110: out_mask = 32'b11111111111111111111111111;
					5'b00111: out_mask = 32'b1111111111111111111111111;
					5'b01000: out_mask = 32'b111111111111111111111111;
					5'b01001: out_mask = 32'b11111111111111111111111;
					5'b01010: out_mask = 32'b1111111111111111111111;
					5'b01011: out_mask = 32'b111111111111111111111;
					5'b01100: out_mask = 32'b11111111111111111111;
					5'b01101: out_mask = 32'b1111111111111111111;
					5'b01110: out_mask = 32'b111111111111111111;
					5'b01111: out_mask = 32'b11111111111111111;
					5'b10000: out_mask = 32'b1111111111111111;
					5'b10001: out_mask = 32'b111111111111111;
					5'b10010: out_mask = 32'b11111111111111;
					5'b10011: out_mask = 32'b1111111111111;
					5'b10100: out_mask = 32'b111111111111;
					5'b10101: out_mask = 32'b11111111111;
					5'b10110: out_mask = 32'b1111111111;
					5'b10111: out_mask = 32'b111111111;
					5'b11000: out_mask = 32'b11111111;
					5'b11001: out_mask = 32'b1111111;
					5'b11010: out_mask = 32'b111111;
					5'b11011: out_mask = 32'b11111;
					5'b11100: out_mask = 32'b1111;
					5'b11101: out_mask = 32'b111;
					5'b11110: out_mask = 32'b11;
					5'b11111: out_mask = 32'b1;
					default: out_mask = 32'b1;
				endcase
			end
			1'b1 : begin  // shift left
				case(in_shift)
					5'b00000: out_mask = 32'b11111111111111111111111111111111;
					5'b00001: out_mask = 32'b11111111111111111111111111111110;
					5'b00010: out_mask = 32'b11111111111111111111111111111100;
					5'b00011: out_mask = 32'b11111111111111111111111111111000;
					5'b00100: out_mask = 32'b11111111111111111111111111110000;
					5'b00101: out_mask = 32'b11111111111111111111111111100000;
					5'b00110: out_mask = 32'b11111111111111111111111111000000;
					5'b00111: out_mask = 32'b11111111111111111111111110000000;
					5'b01000: out_mask = 32'b11111111111111111111111100000000;
					5'b01001: out_mask = 32'b11111111111111111111111000000000;
					5'b01010: out_mask = 32'b11111111111111111111110000000000;
					5'b01011: out_mask = 32'b11111111111111111111100000000000;
					5'b01100: out_mask = 32'b11111111111111111111000000000000;
					5'b01101: out_mask = 32'b11111111111111111110000000000000;
					5'b01110: out_mask = 32'b11111111111111111100000000000000;
					5'b01111: out_mask = 32'b11111111111111111000000000000000;
					5'b10000: out_mask = 32'b11111111111111110000000000000000;
					5'b10001: out_mask = 32'b11111111111111100000000000000000;
					5'b10010: out_mask = 32'b11111111111111000000000000000000;
					5'b10011: out_mask = 32'b11111111111110000000000000000000;
					5'b10100: out_mask = 32'b11111111111100000000000000000000;
					5'b10101: out_mask = 32'b11111111111000000000000000000000;
					5'b10110: out_mask = 32'b11111111110000000000000000000000;
					5'b10111: out_mask = 32'b11111111100000000000000000000000;
					5'b11000: out_mask = 32'b11111111000000000000000000000000;
					5'b11001: out_mask = 32'b11111110000000000000000000000000;
					5'b11010: out_mask = 32'b11111100000000000000000000000000;
					5'b11011: out_mask = 32'b11111000000000000000000000000000;
					5'b11100: out_mask = 32'b11110000000000000000000000000000;
					5'b11101: out_mask = 32'b11100000000000000000000000000000;
					5'b11110: out_mask = 32'b11000000000000000000000000000000;
					5'b11111: out_mask = 32'b10000000000000000000000000000000;
					default: out_mask = 32'b1;
				endcase
			end
			default : out_mask = 32'b1;
		endcase
	end

endmodule

// ----------------------------
